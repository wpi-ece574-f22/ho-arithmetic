module div(input  wire [7:0] y,
	   input wire [7:0]  x,
	   output wire [7:0] r,
	   output wire [7:0] q,
	   input wire 	     start,
	   output wire 	     ready,
	   input wire 	     clk,
	   input wire 	     reset);

   // implement a restoring divider on 8-bit precision
   
endmodule
